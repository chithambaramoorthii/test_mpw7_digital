magic
tech sky130B
magscale 1 2
timestamp 1662565876
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 14 1300 179110 117552
<< metal2 >>
rect 18 119200 74 120000
rect 1306 119200 1362 120000
rect 1950 119200 2006 120000
rect 3238 119200 3294 120000
rect 3882 119200 3938 120000
rect 5170 119200 5226 120000
rect 5814 119200 5870 120000
rect 7102 119200 7158 120000
rect 7746 119200 7802 120000
rect 9034 119200 9090 120000
rect 9678 119200 9734 120000
rect 10966 119200 11022 120000
rect 11610 119200 11666 120000
rect 12898 119200 12954 120000
rect 13542 119200 13598 120000
rect 14830 119200 14886 120000
rect 15474 119200 15530 120000
rect 16762 119200 16818 120000
rect 17406 119200 17462 120000
rect 18694 119200 18750 120000
rect 19338 119200 19394 120000
rect 20626 119200 20682 120000
rect 21270 119200 21326 120000
rect 22558 119200 22614 120000
rect 23202 119200 23258 120000
rect 24490 119200 24546 120000
rect 25134 119200 25190 120000
rect 26422 119200 26478 120000
rect 27066 119200 27122 120000
rect 28354 119200 28410 120000
rect 28998 119200 29054 120000
rect 30286 119200 30342 120000
rect 30930 119200 30986 120000
rect 32218 119200 32274 120000
rect 32862 119200 32918 120000
rect 34150 119200 34206 120000
rect 34794 119200 34850 120000
rect 36082 119200 36138 120000
rect 36726 119200 36782 120000
rect 38014 119200 38070 120000
rect 38658 119200 38714 120000
rect 39946 119200 40002 120000
rect 40590 119200 40646 120000
rect 41878 119200 41934 120000
rect 42522 119200 42578 120000
rect 43810 119200 43866 120000
rect 44454 119200 44510 120000
rect 45742 119200 45798 120000
rect 46386 119200 46442 120000
rect 47674 119200 47730 120000
rect 48318 119200 48374 120000
rect 49606 119200 49662 120000
rect 50250 119200 50306 120000
rect 51538 119200 51594 120000
rect 52182 119200 52238 120000
rect 53470 119200 53526 120000
rect 54758 119200 54814 120000
rect 55402 119200 55458 120000
rect 56690 119200 56746 120000
rect 57334 119200 57390 120000
rect 58622 119200 58678 120000
rect 59266 119200 59322 120000
rect 60554 119200 60610 120000
rect 61198 119200 61254 120000
rect 62486 119200 62542 120000
rect 63130 119200 63186 120000
rect 64418 119200 64474 120000
rect 65062 119200 65118 120000
rect 66350 119200 66406 120000
rect 66994 119200 67050 120000
rect 68282 119200 68338 120000
rect 68926 119200 68982 120000
rect 70214 119200 70270 120000
rect 70858 119200 70914 120000
rect 72146 119200 72202 120000
rect 72790 119200 72846 120000
rect 74078 119200 74134 120000
rect 74722 119200 74778 120000
rect 76010 119200 76066 120000
rect 76654 119200 76710 120000
rect 77942 119200 77998 120000
rect 78586 119200 78642 120000
rect 79874 119200 79930 120000
rect 80518 119200 80574 120000
rect 81806 119200 81862 120000
rect 82450 119200 82506 120000
rect 83738 119200 83794 120000
rect 84382 119200 84438 120000
rect 85670 119200 85726 120000
rect 86314 119200 86370 120000
rect 87602 119200 87658 120000
rect 88246 119200 88302 120000
rect 89534 119200 89590 120000
rect 90178 119200 90234 120000
rect 91466 119200 91522 120000
rect 92110 119200 92166 120000
rect 93398 119200 93454 120000
rect 94042 119200 94098 120000
rect 95330 119200 95386 120000
rect 95974 119200 96030 120000
rect 97262 119200 97318 120000
rect 97906 119200 97962 120000
rect 99194 119200 99250 120000
rect 99838 119200 99894 120000
rect 101126 119200 101182 120000
rect 101770 119200 101826 120000
rect 103058 119200 103114 120000
rect 103702 119200 103758 120000
rect 104990 119200 105046 120000
rect 105634 119200 105690 120000
rect 106922 119200 106978 120000
rect 107566 119200 107622 120000
rect 108854 119200 108910 120000
rect 109498 119200 109554 120000
rect 110786 119200 110842 120000
rect 111430 119200 111486 120000
rect 112718 119200 112774 120000
rect 113362 119200 113418 120000
rect 114650 119200 114706 120000
rect 115294 119200 115350 120000
rect 116582 119200 116638 120000
rect 117226 119200 117282 120000
rect 118514 119200 118570 120000
rect 119158 119200 119214 120000
rect 120446 119200 120502 120000
rect 121090 119200 121146 120000
rect 122378 119200 122434 120000
rect 123022 119200 123078 120000
rect 124310 119200 124366 120000
rect 124954 119200 125010 120000
rect 126242 119200 126298 120000
rect 126886 119200 126942 120000
rect 128174 119200 128230 120000
rect 128818 119200 128874 120000
rect 130106 119200 130162 120000
rect 130750 119200 130806 120000
rect 132038 119200 132094 120000
rect 132682 119200 132738 120000
rect 133970 119200 134026 120000
rect 134614 119200 134670 120000
rect 135902 119200 135958 120000
rect 136546 119200 136602 120000
rect 137834 119200 137890 120000
rect 139122 119200 139178 120000
rect 139766 119200 139822 120000
rect 141054 119200 141110 120000
rect 141698 119200 141754 120000
rect 142986 119200 143042 120000
rect 143630 119200 143686 120000
rect 144918 119200 144974 120000
rect 145562 119200 145618 120000
rect 146850 119200 146906 120000
rect 147494 119200 147550 120000
rect 148782 119200 148838 120000
rect 149426 119200 149482 120000
rect 150714 119200 150770 120000
rect 151358 119200 151414 120000
rect 152646 119200 152702 120000
rect 153290 119200 153346 120000
rect 154578 119200 154634 120000
rect 155222 119200 155278 120000
rect 156510 119200 156566 120000
rect 157154 119200 157210 120000
rect 158442 119200 158498 120000
rect 159086 119200 159142 120000
rect 160374 119200 160430 120000
rect 161018 119200 161074 120000
rect 162306 119200 162362 120000
rect 162950 119200 163006 120000
rect 164238 119200 164294 120000
rect 164882 119200 164938 120000
rect 166170 119200 166226 120000
rect 166814 119200 166870 120000
rect 168102 119200 168158 120000
rect 168746 119200 168802 120000
rect 170034 119200 170090 120000
rect 170678 119200 170734 120000
rect 171966 119200 172022 120000
rect 172610 119200 172666 120000
rect 173898 119200 173954 120000
rect 174542 119200 174598 120000
rect 175830 119200 175886 120000
rect 176474 119200 176530 120000
rect 177762 119200 177818 120000
rect 178406 119200 178462 120000
rect 179694 119200 179750 120000
rect 18 0 74 800
rect 662 0 718 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 50894 0 50950 800
rect 52182 0 52238 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 56690 0 56746 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59910 0 59966 800
rect 60554 0 60610 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63774 0 63830 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 69570 0 69626 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76010 0 76066 800
rect 77298 0 77354 800
rect 77942 0 77998 800
rect 79230 0 79286 800
rect 79874 0 79930 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85026 0 85082 800
rect 86314 0 86370 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 88890 0 88946 800
rect 90178 0 90234 800
rect 90822 0 90878 800
rect 92110 0 92166 800
rect 92754 0 92810 800
rect 94042 0 94098 800
rect 94686 0 94742 800
rect 95974 0 96030 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 98550 0 98606 800
rect 99838 0 99894 800
rect 100482 0 100538 800
rect 101770 0 101826 800
rect 102414 0 102470 800
rect 103702 0 103758 800
rect 104346 0 104402 800
rect 105634 0 105690 800
rect 106278 0 106334 800
rect 107566 0 107622 800
rect 108210 0 108266 800
rect 109498 0 109554 800
rect 110142 0 110198 800
rect 111430 0 111486 800
rect 112074 0 112130 800
rect 113362 0 113418 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 115938 0 115994 800
rect 117226 0 117282 800
rect 117870 0 117926 800
rect 119158 0 119214 800
rect 119802 0 119858 800
rect 121090 0 121146 800
rect 121734 0 121790 800
rect 123022 0 123078 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 125598 0 125654 800
rect 126886 0 126942 800
rect 127530 0 127586 800
rect 128818 0 128874 800
rect 129462 0 129518 800
rect 130750 0 130806 800
rect 131394 0 131450 800
rect 132682 0 132738 800
rect 133326 0 133382 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 136546 0 136602 800
rect 137190 0 137246 800
rect 138478 0 138534 800
rect 139122 0 139178 800
rect 140410 0 140466 800
rect 141054 0 141110 800
rect 142342 0 142398 800
rect 142986 0 143042 800
rect 144274 0 144330 800
rect 144918 0 144974 800
rect 146206 0 146262 800
rect 146850 0 146906 800
rect 148138 0 148194 800
rect 148782 0 148838 800
rect 150070 0 150126 800
rect 150714 0 150770 800
rect 152002 0 152058 800
rect 152646 0 152702 800
rect 153934 0 153990 800
rect 154578 0 154634 800
rect 155866 0 155922 800
rect 156510 0 156566 800
rect 157798 0 157854 800
rect 158442 0 158498 800
rect 159730 0 159786 800
rect 160374 0 160430 800
rect 161662 0 161718 800
rect 162306 0 162362 800
rect 163594 0 163650 800
rect 164238 0 164294 800
rect 165526 0 165582 800
rect 166170 0 166226 800
rect 167458 0 167514 800
rect 168746 0 168802 800
rect 169390 0 169446 800
rect 170678 0 170734 800
rect 171322 0 171378 800
rect 172610 0 172666 800
rect 173254 0 173310 800
rect 174542 0 174598 800
rect 175186 0 175242 800
rect 176474 0 176530 800
rect 177118 0 177174 800
rect 178406 0 178462 800
rect 179050 0 179106 800
<< obsm2 >>
rect 130 119144 1250 119785
rect 1418 119144 1894 119785
rect 2062 119144 3182 119785
rect 3350 119144 3826 119785
rect 3994 119144 5114 119785
rect 5282 119144 5758 119785
rect 5926 119144 7046 119785
rect 7214 119144 7690 119785
rect 7858 119144 8978 119785
rect 9146 119144 9622 119785
rect 9790 119144 10910 119785
rect 11078 119144 11554 119785
rect 11722 119144 12842 119785
rect 13010 119144 13486 119785
rect 13654 119144 14774 119785
rect 14942 119144 15418 119785
rect 15586 119144 16706 119785
rect 16874 119144 17350 119785
rect 17518 119144 18638 119785
rect 18806 119144 19282 119785
rect 19450 119144 20570 119785
rect 20738 119144 21214 119785
rect 21382 119144 22502 119785
rect 22670 119144 23146 119785
rect 23314 119144 24434 119785
rect 24602 119144 25078 119785
rect 25246 119144 26366 119785
rect 26534 119144 27010 119785
rect 27178 119144 28298 119785
rect 28466 119144 28942 119785
rect 29110 119144 30230 119785
rect 30398 119144 30874 119785
rect 31042 119144 32162 119785
rect 32330 119144 32806 119785
rect 32974 119144 34094 119785
rect 34262 119144 34738 119785
rect 34906 119144 36026 119785
rect 36194 119144 36670 119785
rect 36838 119144 37958 119785
rect 38126 119144 38602 119785
rect 38770 119144 39890 119785
rect 40058 119144 40534 119785
rect 40702 119144 41822 119785
rect 41990 119144 42466 119785
rect 42634 119144 43754 119785
rect 43922 119144 44398 119785
rect 44566 119144 45686 119785
rect 45854 119144 46330 119785
rect 46498 119144 47618 119785
rect 47786 119144 48262 119785
rect 48430 119144 49550 119785
rect 49718 119144 50194 119785
rect 50362 119144 51482 119785
rect 51650 119144 52126 119785
rect 52294 119144 53414 119785
rect 53582 119144 54702 119785
rect 54870 119144 55346 119785
rect 55514 119144 56634 119785
rect 56802 119144 57278 119785
rect 57446 119144 58566 119785
rect 58734 119144 59210 119785
rect 59378 119144 60498 119785
rect 60666 119144 61142 119785
rect 61310 119144 62430 119785
rect 62598 119144 63074 119785
rect 63242 119144 64362 119785
rect 64530 119144 65006 119785
rect 65174 119144 66294 119785
rect 66462 119144 66938 119785
rect 67106 119144 68226 119785
rect 68394 119144 68870 119785
rect 69038 119144 70158 119785
rect 70326 119144 70802 119785
rect 70970 119144 72090 119785
rect 72258 119144 72734 119785
rect 72902 119144 74022 119785
rect 74190 119144 74666 119785
rect 74834 119144 75954 119785
rect 76122 119144 76598 119785
rect 76766 119144 77886 119785
rect 78054 119144 78530 119785
rect 78698 119144 79818 119785
rect 79986 119144 80462 119785
rect 80630 119144 81750 119785
rect 81918 119144 82394 119785
rect 82562 119144 83682 119785
rect 83850 119144 84326 119785
rect 84494 119144 85614 119785
rect 85782 119144 86258 119785
rect 86426 119144 87546 119785
rect 87714 119144 88190 119785
rect 88358 119144 89478 119785
rect 89646 119144 90122 119785
rect 90290 119144 91410 119785
rect 91578 119144 92054 119785
rect 92222 119144 93342 119785
rect 93510 119144 93986 119785
rect 94154 119144 95274 119785
rect 95442 119144 95918 119785
rect 96086 119144 97206 119785
rect 97374 119144 97850 119785
rect 98018 119144 99138 119785
rect 99306 119144 99782 119785
rect 99950 119144 101070 119785
rect 101238 119144 101714 119785
rect 101882 119144 103002 119785
rect 103170 119144 103646 119785
rect 103814 119144 104934 119785
rect 105102 119144 105578 119785
rect 105746 119144 106866 119785
rect 107034 119144 107510 119785
rect 107678 119144 108798 119785
rect 108966 119144 109442 119785
rect 109610 119144 110730 119785
rect 110898 119144 111374 119785
rect 111542 119144 112662 119785
rect 112830 119144 113306 119785
rect 113474 119144 114594 119785
rect 114762 119144 115238 119785
rect 115406 119144 116526 119785
rect 116694 119144 117170 119785
rect 117338 119144 118458 119785
rect 118626 119144 119102 119785
rect 119270 119144 120390 119785
rect 120558 119144 121034 119785
rect 121202 119144 122322 119785
rect 122490 119144 122966 119785
rect 123134 119144 124254 119785
rect 124422 119144 124898 119785
rect 125066 119144 126186 119785
rect 126354 119144 126830 119785
rect 126998 119144 128118 119785
rect 128286 119144 128762 119785
rect 128930 119144 130050 119785
rect 130218 119144 130694 119785
rect 130862 119144 131982 119785
rect 132150 119144 132626 119785
rect 132794 119144 133914 119785
rect 134082 119144 134558 119785
rect 134726 119144 135846 119785
rect 136014 119144 136490 119785
rect 136658 119144 137778 119785
rect 137946 119144 139066 119785
rect 139234 119144 139710 119785
rect 139878 119144 140998 119785
rect 141166 119144 141642 119785
rect 141810 119144 142930 119785
rect 143098 119144 143574 119785
rect 143742 119144 144862 119785
rect 145030 119144 145506 119785
rect 145674 119144 146794 119785
rect 146962 119144 147438 119785
rect 147606 119144 148726 119785
rect 148894 119144 149370 119785
rect 149538 119144 150658 119785
rect 150826 119144 151302 119785
rect 151470 119144 152590 119785
rect 152758 119144 153234 119785
rect 153402 119144 154522 119785
rect 154690 119144 155166 119785
rect 155334 119144 156454 119785
rect 156622 119144 157098 119785
rect 157266 119144 158386 119785
rect 158554 119144 159030 119785
rect 159198 119144 160318 119785
rect 160486 119144 160962 119785
rect 161130 119144 162250 119785
rect 162418 119144 162894 119785
rect 163062 119144 164182 119785
rect 164350 119144 164826 119785
rect 164994 119144 166114 119785
rect 166282 119144 166758 119785
rect 166926 119144 168046 119785
rect 168214 119144 168690 119785
rect 168858 119144 169978 119785
rect 170146 119144 170622 119785
rect 170790 119144 171910 119785
rect 172078 119144 172554 119785
rect 172722 119144 173842 119785
rect 174010 119144 174486 119785
rect 174654 119144 175774 119785
rect 175942 119144 176418 119785
rect 176586 119144 177706 119785
rect 177874 119144 178350 119785
rect 178518 119144 179104 119785
rect 20 856 179104 119144
rect 130 31 606 856
rect 774 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7690 856
rect 7858 31 8334 856
rect 8502 31 9622 856
rect 9790 31 10266 856
rect 10434 31 11554 856
rect 11722 31 12198 856
rect 12366 31 13486 856
rect 13654 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16062 856
rect 16230 31 17350 856
rect 17518 31 17994 856
rect 18162 31 19282 856
rect 19450 31 19926 856
rect 20094 31 21214 856
rect 21382 31 21858 856
rect 22026 31 23146 856
rect 23314 31 23790 856
rect 23958 31 25078 856
rect 25246 31 25722 856
rect 25890 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28942 856
rect 29110 31 29586 856
rect 29754 31 30874 856
rect 31042 31 31518 856
rect 31686 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36670 856
rect 36838 31 37314 856
rect 37482 31 38602 856
rect 38770 31 39246 856
rect 39414 31 40534 856
rect 40702 31 41178 856
rect 41346 31 42466 856
rect 42634 31 43110 856
rect 43278 31 44398 856
rect 44566 31 45042 856
rect 45210 31 46330 856
rect 46498 31 46974 856
rect 47142 31 48262 856
rect 48430 31 48906 856
rect 49074 31 50194 856
rect 50362 31 50838 856
rect 51006 31 52126 856
rect 52294 31 52770 856
rect 52938 31 54058 856
rect 54226 31 54702 856
rect 54870 31 55990 856
rect 56158 31 56634 856
rect 56802 31 57922 856
rect 58090 31 58566 856
rect 58734 31 59854 856
rect 60022 31 60498 856
rect 60666 31 61786 856
rect 61954 31 62430 856
rect 62598 31 63718 856
rect 63886 31 64362 856
rect 64530 31 65650 856
rect 65818 31 66294 856
rect 66462 31 67582 856
rect 67750 31 68226 856
rect 68394 31 69514 856
rect 69682 31 70158 856
rect 70326 31 71446 856
rect 71614 31 72090 856
rect 72258 31 73378 856
rect 73546 31 74022 856
rect 74190 31 75310 856
rect 75478 31 75954 856
rect 76122 31 77242 856
rect 77410 31 77886 856
rect 78054 31 79174 856
rect 79342 31 79818 856
rect 79986 31 81106 856
rect 81274 31 81750 856
rect 81918 31 83038 856
rect 83206 31 84326 856
rect 84494 31 84970 856
rect 85138 31 86258 856
rect 86426 31 86902 856
rect 87070 31 88190 856
rect 88358 31 88834 856
rect 89002 31 90122 856
rect 90290 31 90766 856
rect 90934 31 92054 856
rect 92222 31 92698 856
rect 92866 31 93986 856
rect 94154 31 94630 856
rect 94798 31 95918 856
rect 96086 31 96562 856
rect 96730 31 97850 856
rect 98018 31 98494 856
rect 98662 31 99782 856
rect 99950 31 100426 856
rect 100594 31 101714 856
rect 101882 31 102358 856
rect 102526 31 103646 856
rect 103814 31 104290 856
rect 104458 31 105578 856
rect 105746 31 106222 856
rect 106390 31 107510 856
rect 107678 31 108154 856
rect 108322 31 109442 856
rect 109610 31 110086 856
rect 110254 31 111374 856
rect 111542 31 112018 856
rect 112186 31 113306 856
rect 113474 31 113950 856
rect 114118 31 115238 856
rect 115406 31 115882 856
rect 116050 31 117170 856
rect 117338 31 117814 856
rect 117982 31 119102 856
rect 119270 31 119746 856
rect 119914 31 121034 856
rect 121202 31 121678 856
rect 121846 31 122966 856
rect 123134 31 123610 856
rect 123778 31 124898 856
rect 125066 31 125542 856
rect 125710 31 126830 856
rect 126998 31 127474 856
rect 127642 31 128762 856
rect 128930 31 129406 856
rect 129574 31 130694 856
rect 130862 31 131338 856
rect 131506 31 132626 856
rect 132794 31 133270 856
rect 133438 31 134558 856
rect 134726 31 135202 856
rect 135370 31 136490 856
rect 136658 31 137134 856
rect 137302 31 138422 856
rect 138590 31 139066 856
rect 139234 31 140354 856
rect 140522 31 140998 856
rect 141166 31 142286 856
rect 142454 31 142930 856
rect 143098 31 144218 856
rect 144386 31 144862 856
rect 145030 31 146150 856
rect 146318 31 146794 856
rect 146962 31 148082 856
rect 148250 31 148726 856
rect 148894 31 150014 856
rect 150182 31 150658 856
rect 150826 31 151946 856
rect 152114 31 152590 856
rect 152758 31 153878 856
rect 154046 31 154522 856
rect 154690 31 155810 856
rect 155978 31 156454 856
rect 156622 31 157742 856
rect 157910 31 158386 856
rect 158554 31 159674 856
rect 159842 31 160318 856
rect 160486 31 161606 856
rect 161774 31 162250 856
rect 162418 31 163538 856
rect 163706 31 164182 856
rect 164350 31 165470 856
rect 165638 31 166114 856
rect 166282 31 167402 856
rect 167570 31 168690 856
rect 168858 31 169334 856
rect 169502 31 170622 856
rect 170790 31 171266 856
rect 171434 31 172554 856
rect 172722 31 173198 856
rect 173366 31 174486 856
rect 174654 31 175130 856
rect 175298 31 176418 856
rect 176586 31 177062 856
rect 177230 31 178350 856
rect 178518 31 178994 856
<< metal3 >>
rect 0 119688 800 119808
rect 179200 119688 180000 119808
rect 0 118328 800 118448
rect 179200 118328 180000 118448
rect 0 117648 800 117768
rect 179200 117648 180000 117768
rect 0 116288 800 116408
rect 179200 116288 180000 116408
rect 0 115608 800 115728
rect 179200 115608 180000 115728
rect 0 114248 800 114368
rect 179200 114248 180000 114368
rect 0 113568 800 113688
rect 179200 113568 180000 113688
rect 0 112208 800 112328
rect 179200 112208 180000 112328
rect 0 111528 800 111648
rect 179200 111528 180000 111648
rect 0 110168 800 110288
rect 179200 110168 180000 110288
rect 0 109488 800 109608
rect 179200 109488 180000 109608
rect 0 108128 800 108248
rect 179200 108128 180000 108248
rect 0 107448 800 107568
rect 179200 107448 180000 107568
rect 0 106088 800 106208
rect 179200 106088 180000 106208
rect 0 105408 800 105528
rect 179200 105408 180000 105528
rect 0 104048 800 104168
rect 179200 104048 180000 104168
rect 0 103368 800 103488
rect 179200 103368 180000 103488
rect 0 102008 800 102128
rect 179200 102008 180000 102128
rect 0 101328 800 101448
rect 179200 101328 180000 101448
rect 0 99968 800 100088
rect 179200 99968 180000 100088
rect 0 99288 800 99408
rect 179200 99288 180000 99408
rect 0 97928 800 98048
rect 179200 97928 180000 98048
rect 0 97248 800 97368
rect 179200 97248 180000 97368
rect 0 95888 800 96008
rect 179200 95888 180000 96008
rect 0 95208 800 95328
rect 179200 95208 180000 95328
rect 0 93848 800 93968
rect 179200 93848 180000 93968
rect 0 93168 800 93288
rect 179200 93168 180000 93288
rect 0 91808 800 91928
rect 179200 91808 180000 91928
rect 0 91128 800 91248
rect 179200 91128 180000 91248
rect 0 89768 800 89888
rect 179200 89768 180000 89888
rect 0 89088 800 89208
rect 179200 89088 180000 89208
rect 0 87728 800 87848
rect 179200 87728 180000 87848
rect 179200 87048 180000 87168
rect 0 86368 800 86488
rect 0 85688 800 85808
rect 179200 85688 180000 85808
rect 179200 85008 180000 85128
rect 0 84328 800 84448
rect 0 83648 800 83768
rect 179200 83648 180000 83768
rect 179200 82968 180000 83088
rect 0 82288 800 82408
rect 0 81608 800 81728
rect 179200 81608 180000 81728
rect 179200 80928 180000 81048
rect 0 80248 800 80368
rect 0 79568 800 79688
rect 179200 79568 180000 79688
rect 179200 78888 180000 79008
rect 0 78208 800 78328
rect 0 77528 800 77648
rect 179200 77528 180000 77648
rect 179200 76848 180000 76968
rect 0 76168 800 76288
rect 0 75488 800 75608
rect 179200 75488 180000 75608
rect 0 74128 800 74248
rect 179200 74128 180000 74248
rect 0 73448 800 73568
rect 179200 73448 180000 73568
rect 0 72088 800 72208
rect 179200 72088 180000 72208
rect 0 71408 800 71528
rect 179200 71408 180000 71528
rect 0 70048 800 70168
rect 179200 70048 180000 70168
rect 0 69368 800 69488
rect 179200 69368 180000 69488
rect 0 68008 800 68128
rect 179200 68008 180000 68128
rect 0 67328 800 67448
rect 179200 67328 180000 67448
rect 0 65968 800 66088
rect 179200 65968 180000 66088
rect 0 65288 800 65408
rect 179200 65288 180000 65408
rect 0 63928 800 64048
rect 179200 63928 180000 64048
rect 0 63248 800 63368
rect 179200 63248 180000 63368
rect 0 61888 800 62008
rect 179200 61888 180000 62008
rect 0 61208 800 61328
rect 179200 61208 180000 61328
rect 0 59848 800 59968
rect 179200 59848 180000 59968
rect 0 59168 800 59288
rect 179200 59168 180000 59288
rect 0 57808 800 57928
rect 179200 57808 180000 57928
rect 0 57128 800 57248
rect 179200 57128 180000 57248
rect 0 55768 800 55888
rect 179200 55768 180000 55888
rect 0 55088 800 55208
rect 179200 55088 180000 55208
rect 0 53728 800 53848
rect 179200 53728 180000 53848
rect 0 53048 800 53168
rect 179200 53048 180000 53168
rect 0 51688 800 51808
rect 179200 51688 180000 51808
rect 0 51008 800 51128
rect 179200 51008 180000 51128
rect 0 49648 800 49768
rect 179200 49648 180000 49768
rect 0 48968 800 49088
rect 179200 48968 180000 49088
rect 0 47608 800 47728
rect 179200 47608 180000 47728
rect 0 46928 800 47048
rect 179200 46928 180000 47048
rect 0 45568 800 45688
rect 179200 45568 180000 45688
rect 0 44888 800 45008
rect 179200 44888 180000 45008
rect 0 43528 800 43648
rect 179200 43528 180000 43648
rect 0 42848 800 42968
rect 179200 42848 180000 42968
rect 0 41488 800 41608
rect 179200 41488 180000 41608
rect 0 40808 800 40928
rect 179200 40808 180000 40928
rect 0 39448 800 39568
rect 179200 39448 180000 39568
rect 0 38768 800 38888
rect 179200 38768 180000 38888
rect 0 37408 800 37528
rect 179200 37408 180000 37528
rect 0 36728 800 36848
rect 179200 36728 180000 36848
rect 0 35368 800 35488
rect 179200 35368 180000 35488
rect 0 34688 800 34808
rect 179200 34688 180000 34808
rect 0 33328 800 33448
rect 179200 33328 180000 33448
rect 0 32648 800 32768
rect 179200 32648 180000 32768
rect 0 31288 800 31408
rect 179200 31288 180000 31408
rect 0 30608 800 30728
rect 179200 30608 180000 30728
rect 0 29248 800 29368
rect 179200 29248 180000 29368
rect 0 28568 800 28688
rect 179200 28568 180000 28688
rect 0 27208 800 27328
rect 179200 27208 180000 27328
rect 0 26528 800 26648
rect 179200 26528 180000 26648
rect 0 25168 800 25288
rect 179200 25168 180000 25288
rect 0 24488 800 24608
rect 179200 24488 180000 24608
rect 0 23128 800 23248
rect 179200 23128 180000 23248
rect 0 22448 800 22568
rect 179200 22448 180000 22568
rect 0 21088 800 21208
rect 179200 21088 180000 21208
rect 0 20408 800 20528
rect 179200 20408 180000 20528
rect 0 19048 800 19168
rect 179200 19048 180000 19168
rect 0 18368 800 18488
rect 179200 18368 180000 18488
rect 0 17008 800 17128
rect 179200 17008 180000 17128
rect 0 16328 800 16448
rect 179200 16328 180000 16448
rect 0 14968 800 15088
rect 179200 14968 180000 15088
rect 0 14288 800 14408
rect 179200 14288 180000 14408
rect 0 12928 800 13048
rect 179200 12928 180000 13048
rect 0 12248 800 12368
rect 179200 12248 180000 12368
rect 0 10888 800 11008
rect 179200 10888 180000 11008
rect 0 10208 800 10328
rect 179200 10208 180000 10328
rect 0 8848 800 8968
rect 179200 8848 180000 8968
rect 0 8168 800 8288
rect 179200 8168 180000 8288
rect 0 6808 800 6928
rect 179200 6808 180000 6928
rect 0 6128 800 6248
rect 179200 6128 180000 6248
rect 0 4768 800 4888
rect 179200 4768 180000 4888
rect 0 4088 800 4208
rect 179200 4088 180000 4208
rect 0 2728 800 2848
rect 179200 2728 180000 2848
rect 0 2048 800 2168
rect 179200 2048 180000 2168
rect 0 688 800 808
rect 179200 688 180000 808
rect 179200 8 180000 128
<< obsm3 >>
rect 880 119608 179120 119781
rect 800 118528 179200 119608
rect 880 118248 179120 118528
rect 800 117848 179200 118248
rect 880 117568 179120 117848
rect 800 116488 179200 117568
rect 880 116208 179120 116488
rect 800 115808 179200 116208
rect 880 115528 179120 115808
rect 800 114448 179200 115528
rect 880 114168 179120 114448
rect 800 113768 179200 114168
rect 880 113488 179120 113768
rect 800 112408 179200 113488
rect 880 112128 179120 112408
rect 800 111728 179200 112128
rect 880 111448 179120 111728
rect 800 110368 179200 111448
rect 880 110088 179120 110368
rect 800 109688 179200 110088
rect 880 109408 179120 109688
rect 800 108328 179200 109408
rect 880 108048 179120 108328
rect 800 107648 179200 108048
rect 880 107368 179120 107648
rect 800 106288 179200 107368
rect 880 106008 179120 106288
rect 800 105608 179200 106008
rect 880 105328 179120 105608
rect 800 104248 179200 105328
rect 880 103968 179120 104248
rect 800 103568 179200 103968
rect 880 103288 179120 103568
rect 800 102208 179200 103288
rect 880 101928 179120 102208
rect 800 101528 179200 101928
rect 880 101248 179120 101528
rect 800 100168 179200 101248
rect 880 99888 179120 100168
rect 800 99488 179200 99888
rect 880 99208 179120 99488
rect 800 98128 179200 99208
rect 880 97848 179120 98128
rect 800 97448 179200 97848
rect 880 97168 179120 97448
rect 800 96088 179200 97168
rect 880 95808 179120 96088
rect 800 95408 179200 95808
rect 880 95128 179120 95408
rect 800 94048 179200 95128
rect 880 93768 179120 94048
rect 800 93368 179200 93768
rect 880 93088 179120 93368
rect 800 92008 179200 93088
rect 880 91728 179120 92008
rect 800 91328 179200 91728
rect 880 91048 179120 91328
rect 800 89968 179200 91048
rect 880 89688 179120 89968
rect 800 89288 179200 89688
rect 880 89008 179120 89288
rect 800 87928 179200 89008
rect 880 87648 179120 87928
rect 800 87248 179200 87648
rect 800 86968 179120 87248
rect 800 86568 179200 86968
rect 880 86288 179200 86568
rect 800 85888 179200 86288
rect 880 85608 179120 85888
rect 800 85208 179200 85608
rect 800 84928 179120 85208
rect 800 84528 179200 84928
rect 880 84248 179200 84528
rect 800 83848 179200 84248
rect 880 83568 179120 83848
rect 800 83168 179200 83568
rect 800 82888 179120 83168
rect 800 82488 179200 82888
rect 880 82208 179200 82488
rect 800 81808 179200 82208
rect 880 81528 179120 81808
rect 800 81128 179200 81528
rect 800 80848 179120 81128
rect 800 80448 179200 80848
rect 880 80168 179200 80448
rect 800 79768 179200 80168
rect 880 79488 179120 79768
rect 800 79088 179200 79488
rect 800 78808 179120 79088
rect 800 78408 179200 78808
rect 880 78128 179200 78408
rect 800 77728 179200 78128
rect 880 77448 179120 77728
rect 800 77048 179200 77448
rect 800 76768 179120 77048
rect 800 76368 179200 76768
rect 880 76088 179200 76368
rect 800 75688 179200 76088
rect 880 75408 179120 75688
rect 800 74328 179200 75408
rect 880 74048 179120 74328
rect 800 73648 179200 74048
rect 880 73368 179120 73648
rect 800 72288 179200 73368
rect 880 72008 179120 72288
rect 800 71608 179200 72008
rect 880 71328 179120 71608
rect 800 70248 179200 71328
rect 880 69968 179120 70248
rect 800 69568 179200 69968
rect 880 69288 179120 69568
rect 800 68208 179200 69288
rect 880 67928 179120 68208
rect 800 67528 179200 67928
rect 880 67248 179120 67528
rect 800 66168 179200 67248
rect 880 65888 179120 66168
rect 800 65488 179200 65888
rect 880 65208 179120 65488
rect 800 64128 179200 65208
rect 880 63848 179120 64128
rect 800 63448 179200 63848
rect 880 63168 179120 63448
rect 800 62088 179200 63168
rect 880 61808 179120 62088
rect 800 61408 179200 61808
rect 880 61128 179120 61408
rect 800 60048 179200 61128
rect 880 59768 179120 60048
rect 800 59368 179200 59768
rect 880 59088 179120 59368
rect 800 58008 179200 59088
rect 880 57728 179120 58008
rect 800 57328 179200 57728
rect 880 57048 179120 57328
rect 800 55968 179200 57048
rect 880 55688 179120 55968
rect 800 55288 179200 55688
rect 880 55008 179120 55288
rect 800 53928 179200 55008
rect 880 53648 179120 53928
rect 800 53248 179200 53648
rect 880 52968 179120 53248
rect 800 51888 179200 52968
rect 880 51608 179120 51888
rect 800 51208 179200 51608
rect 880 50928 179120 51208
rect 800 49848 179200 50928
rect 880 49568 179120 49848
rect 800 49168 179200 49568
rect 880 48888 179120 49168
rect 800 47808 179200 48888
rect 880 47528 179120 47808
rect 800 47128 179200 47528
rect 880 46848 179120 47128
rect 800 45768 179200 46848
rect 880 45488 179120 45768
rect 800 45088 179200 45488
rect 880 44808 179120 45088
rect 800 43728 179200 44808
rect 880 43448 179120 43728
rect 800 43048 179200 43448
rect 880 42768 179120 43048
rect 800 41688 179200 42768
rect 880 41408 179120 41688
rect 800 41008 179200 41408
rect 880 40728 179120 41008
rect 800 39648 179200 40728
rect 880 39368 179120 39648
rect 800 38968 179200 39368
rect 880 38688 179120 38968
rect 800 37608 179200 38688
rect 880 37328 179120 37608
rect 800 36928 179200 37328
rect 880 36648 179120 36928
rect 800 35568 179200 36648
rect 880 35288 179120 35568
rect 800 34888 179200 35288
rect 880 34608 179120 34888
rect 800 33528 179200 34608
rect 880 33248 179120 33528
rect 800 32848 179200 33248
rect 880 32568 179120 32848
rect 800 31488 179200 32568
rect 880 31208 179120 31488
rect 800 30808 179200 31208
rect 880 30528 179120 30808
rect 800 29448 179200 30528
rect 880 29168 179120 29448
rect 800 28768 179200 29168
rect 880 28488 179120 28768
rect 800 27408 179200 28488
rect 880 27128 179120 27408
rect 800 26728 179200 27128
rect 880 26448 179120 26728
rect 800 25368 179200 26448
rect 880 25088 179120 25368
rect 800 24688 179200 25088
rect 880 24408 179120 24688
rect 800 23328 179200 24408
rect 880 23048 179120 23328
rect 800 22648 179200 23048
rect 880 22368 179120 22648
rect 800 21288 179200 22368
rect 880 21008 179120 21288
rect 800 20608 179200 21008
rect 880 20328 179120 20608
rect 800 19248 179200 20328
rect 880 18968 179120 19248
rect 800 18568 179200 18968
rect 880 18288 179120 18568
rect 800 17208 179200 18288
rect 880 16928 179120 17208
rect 800 16528 179200 16928
rect 880 16248 179120 16528
rect 800 15168 179200 16248
rect 880 14888 179120 15168
rect 800 14488 179200 14888
rect 880 14208 179120 14488
rect 800 13128 179200 14208
rect 880 12848 179120 13128
rect 800 12448 179200 12848
rect 880 12168 179120 12448
rect 800 11088 179200 12168
rect 880 10808 179120 11088
rect 800 10408 179200 10808
rect 880 10128 179120 10408
rect 800 9048 179200 10128
rect 880 8768 179120 9048
rect 800 8368 179200 8768
rect 880 8088 179120 8368
rect 800 7008 179200 8088
rect 880 6728 179120 7008
rect 800 6328 179200 6728
rect 880 6048 179120 6328
rect 800 4968 179200 6048
rect 880 4688 179120 4968
rect 800 4288 179200 4688
rect 880 4008 179120 4288
rect 800 2928 179200 4008
rect 880 2648 179120 2928
rect 800 2248 179200 2648
rect 880 1968 179120 2248
rect 800 888 179200 1968
rect 880 608 179120 888
rect 800 208 179200 608
rect 800 35 179120 208
<< metal4 >>
rect 4208 2128 4528 117552
rect 9316 17360 9636 32688
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 40355 20163 40421 106861
<< labels >>
rlabel metal2 s 144274 0 144330 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 179200 34688 180000 34808 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 80518 119200 80574 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 179200 67328 180000 67448 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 72790 119200 72846 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 179200 113568 180000 113688 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 85670 119200 85726 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 68282 119200 68338 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 76010 119200 76066 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 179200 80928 180000 81048 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 36082 119200 36138 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 124310 119200 124366 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 70858 119200 70914 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 97906 119200 97962 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5814 119200 5870 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 132038 119200 132094 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 117226 119200 117282 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 179200 68008 180000 68128 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 171966 119200 172022 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 179200 57128 180000 57248 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 101770 119200 101826 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 179200 21088 180000 21208 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 179200 18368 180000 18488 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 119158 119200 119214 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 82450 119200 82506 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 56690 119200 56746 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 179200 22448 180000 22568 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 30930 119200 30986 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 34150 119200 34206 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 57334 119200 57390 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 132682 119200 132738 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 179200 29248 180000 29368 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 179200 118328 180000 118448 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 18 119200 74 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 47674 119200 47730 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 121090 119200 121146 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 179200 79568 180000 79688 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 179200 99288 180000 99408 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 14830 119200 14886 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 49606 119200 49662 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 36726 119200 36782 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 58622 119200 58678 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 144918 119200 144974 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 137834 119200 137890 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 174542 119200 174598 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 45742 119200 45798 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 170678 119200 170734 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 179200 109488 180000 109608 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 179200 85688 180000 85808 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 179200 2048 180000 2168 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 179200 65968 180000 66088 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 179200 104048 180000 104168 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 179200 87048 180000 87168 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 27066 119200 27122 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 140410 0 140466 800 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 60554 119200 60610 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 179200 51688 180000 51808 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 173898 119200 173954 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 179200 102008 180000 102128 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 179200 82968 180000 83088 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 178406 119200 178462 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 179200 70048 180000 70168 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 59266 119200 59322 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 179200 61888 180000 62008 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 105634 119200 105690 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 91466 119200 91522 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 28354 119200 28410 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 179200 28568 180000 28688 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 148782 119200 148838 120000 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 179200 44888 180000 45008 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 179200 10208 180000 10328 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 95974 119200 96030 120000 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 54758 119200 54814 120000 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 179200 107448 180000 107568 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 179200 63248 180000 63368 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 111430 119200 111486 120000 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 179200 6808 180000 6928 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 136546 119200 136602 120000 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 179200 63928 180000 64048 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 1306 119200 1362 120000 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 141054 119200 141110 120000 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 90178 119200 90234 120000 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 150714 119200 150770 120000 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 179200 59168 180000 59288 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 130750 119200 130806 120000 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 38014 119200 38070 120000 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 179200 77528 180000 77648 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 179200 31288 180000 31408 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 179200 95888 180000 96008 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 143630 119200 143686 120000 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 32862 119200 32918 120000 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 179200 47608 180000 47728 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 179200 89768 180000 89888 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 179200 57808 180000 57928 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 84382 119200 84438 120000 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 99194 119200 99250 120000 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 7746 119200 7802 120000 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 147494 119200 147550 120000 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 175830 119200 175886 120000 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 179200 33328 180000 33448 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 179200 36728 180000 36848 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 179200 85008 180000 85128 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 79874 119200 79930 120000 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 135902 119200 135958 120000 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 32218 119200 32274 120000 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 172610 119200 172666 120000 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 662 0 718 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 154578 119200 154634 120000 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 41878 119200 41934 120000 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 179200 4088 180000 4208 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 179200 111528 180000 111648 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 23202 119200 23258 120000 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 92110 119200 92166 120000 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 179200 78888 180000 79008 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 179200 27208 180000 27328 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 179200 4768 180000 4888 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 66994 119200 67050 120000 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 179200 65288 180000 65408 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 179200 89088 180000 89208 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 179200 8848 180000 8968 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 179200 14288 180000 14408 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 179200 14968 180000 15088 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 155222 119200 155278 120000 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 688 800 808 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 89534 119200 89590 120000 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 179200 75488 180000 75608 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 81806 119200 81862 120000 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 65062 119200 65118 120000 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 116582 119200 116638 120000 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 34794 119200 34850 120000 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 13542 119200 13598 120000 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 179200 38768 180000 38888 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 168746 119200 168802 120000 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 12898 119200 12954 120000 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 179200 23128 180000 23248 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 179200 49648 180000 49768 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 64418 119200 64474 120000 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 1950 119200 2006 120000 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 107566 119200 107622 120000 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 120446 119200 120502 120000 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 139766 119200 139822 120000 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 166170 119200 166226 120000 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 93398 119200 93454 120000 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 179200 101328 180000 101448 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 179200 688 180000 808 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 55402 119200 55458 120000 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 168102 119200 168158 120000 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 3238 119200 3294 120000 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 179200 103368 180000 103488 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 179200 35368 180000 35488 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 179200 42848 180000 42968 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 42522 119200 42578 120000 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 40590 119200 40646 120000 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 179200 115608 180000 115728 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 128174 119200 128230 120000 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 179200 24488 180000 24608 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 113362 119200 113418 120000 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 179200 37408 180000 37528 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 21270 119200 21326 120000 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 62486 119200 62542 120000 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 162306 119200 162362 120000 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 149426 119200 149482 120000 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 179200 8168 180000 8288 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 87602 119200 87658 120000 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 76654 119200 76710 120000 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 72146 119200 72202 120000 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 177762 119200 177818 120000 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 83738 119200 83794 120000 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 179200 43528 180000 43648 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 179200 39448 180000 39568 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 170034 119200 170090 120000 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 145562 119200 145618 120000 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 103058 119200 103114 120000 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 10966 119200 11022 120000 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 179200 48968 180000 49088 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 179200 8 180000 128 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 164882 119200 164938 120000 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 88246 119200 88302 120000 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 24490 119200 24546 120000 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 104990 119200 105046 120000 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 20626 119200 20682 120000 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 63130 119200 63186 120000 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 52182 119200 52238 120000 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 179200 45568 180000 45688 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 112718 119200 112774 120000 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 108854 119200 108910 120000 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 109498 119200 109554 120000 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 157154 119200 157210 120000 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 78586 119200 78642 120000 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 94042 119200 94098 120000 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 44454 119200 44510 120000 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 153290 119200 153346 120000 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 179200 117648 180000 117768 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 9034 119200 9090 120000 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 156510 119200 156566 120000 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 179200 55088 180000 55208 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 99838 119200 99894 120000 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 176474 119200 176530 120000 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 179200 53048 180000 53168 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 128818 119200 128874 120000 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 146850 119200 146906 120000 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 179200 83648 180000 83768 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 118514 119200 118570 120000 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 179200 112208 180000 112328 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 179200 26528 180000 26648 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 179200 53728 180000 53848 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 179200 93848 180000 93968 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 179200 6128 180000 6248 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 179200 72088 180000 72208 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 179200 110168 180000 110288 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 179200 30608 180000 30728 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 161018 119200 161074 120000 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 179200 51008 180000 51128 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 179694 119200 179750 120000 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 162950 119200 163006 120000 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 74078 119200 74134 120000 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 48318 119200 48374 120000 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 179200 16328 180000 16448 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 179200 55768 180000 55888 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 179200 91808 180000 91928 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 166814 119200 166870 120000 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 11610 119200 11666 120000 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 38658 119200 38714 120000 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 179200 12928 180000 13048 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 179200 93168 180000 93288 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 101126 119200 101182 120000 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 77942 119200 77998 120000 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 179200 108128 180000 108248 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 68926 119200 68982 120000 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 179200 91128 180000 91248 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 134614 119200 134670 120000 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 22558 119200 22614 120000 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 151358 119200 151414 120000 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 159086 119200 159142 120000 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 160374 119200 160430 120000 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 110786 119200 110842 120000 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 26422 119200 26478 120000 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 106922 119200 106978 120000 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 179200 73448 180000 73568 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 179200 106088 180000 106208 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 179200 97928 180000 98048 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 86314 119200 86370 120000 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 179200 76848 180000 76968 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 179200 2728 180000 2848 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 74722 119200 74778 120000 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 18694 119200 18750 120000 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 179200 97248 180000 97368 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 30286 119200 30342 120000 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 123022 119200 123078 120000 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 25134 119200 25190 120000 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 39946 119200 40002 120000 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 9316 17360 9636 32688 6 vssd1
port 503 nsew ground bidirectional
rlabel metal3 s 179200 12248 180000 12368 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 16762 119200 16818 120000 6 wb_rst_i
port 505 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 95330 119200 95386 120000 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 61198 119200 61254 120000 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal3 s 179200 105408 180000 105528 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal3 s 179200 95208 180000 95328 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal3 s 179200 32648 180000 32768 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 97262 119200 97318 120000 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 142986 119200 143042 120000 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal3 s 179200 17008 180000 17128 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 15474 119200 15530 120000 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 51538 119200 51594 120000 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal3 s 179200 74128 180000 74248 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 164238 119200 164294 120000 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 124954 119200 125010 120000 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal3 s 179200 46928 180000 47048 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 122378 119200 122434 120000 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal3 s 179200 20408 180000 20528 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 53470 119200 53526 120000 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal3 s 179200 119688 180000 119808 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal3 s 179200 59848 180000 59968 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 114650 119200 114706 120000 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 152646 119200 152702 120000 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 17406 119200 17462 120000 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal3 s 179200 71408 180000 71528 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 158442 119200 158498 120000 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal3 s 179200 99968 180000 100088 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal3 s 179200 25168 180000 25288 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 141698 119200 141754 120000 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 50250 119200 50306 120000 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal3 s 179200 69368 180000 69488 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal3 s 179200 19048 180000 19168 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal3 s 179200 40808 180000 40928 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 139122 119200 139178 120000 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal3 s 179200 114248 180000 114368 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal3 s 179200 61208 180000 61328 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal3 s 179200 116288 180000 116408 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 133970 119200 134026 120000 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 168746 0 168802 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 66350 119200 66406 120000 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 103702 119200 103758 120000 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 70214 119200 70270 120000 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 130106 119200 130162 120000 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal3 s 179200 10888 180000 11008 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal3 s 179200 87728 180000 87848 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal3 s 179200 81608 180000 81728 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 126886 119200 126942 120000 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 126242 119200 126298 120000 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 19338 119200 19394 120000 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 46386 119200 46442 120000 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 7102 119200 7158 120000 6 wbs_stb_i
port 608 nsew signal input
rlabel metal3 s 179200 41488 180000 41608 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7851504
string GDS_FILE /home/nvm_user4/usr/mpw_7_files/caravel_user_project/openlane/user_proj_example/runs/22_09_07_21_19/results/signoff/user_proj_example.magic.gds
string GDS_START 404892
<< end >>

